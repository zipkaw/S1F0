module cpu #(
    parameters
) (
    ports
);
    
endmodule